let's start boizzzz